module inst

pub enum Opcode {
	hlt
	ldc
	add
	sub
	mul
	div
	jmp
	jmpf
	jmpb
}
