module inst

pub enum Opcode {
	hlt
	ldc
	add
	sub
	mul
	div
	inc
	dec
	jmp
	jeq
	jmpf
	jmpb
	eq
	neq
	gt
	gte
	lt
	lte
	inv
}
