module inst

pub struct Instruction {
	opcode Opcode
}
