module test

import @asm { Visitor }
import inst { Instruction }
import vm
