module test
import @asm
import inst
import vm

