module inst

pub struct Instruction {
pub:
	opcode Opcode
	bits   []int
}
