module inst

pub enum Opcode {
	hlt
}
